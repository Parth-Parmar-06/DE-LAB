module not_2(output Y, input A);
	not(Y,A);
endmodule