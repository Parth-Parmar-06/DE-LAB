module or_2(output Y, input A,B);
	or(Y,A,B);
endmodule