module and_1(output Y, input A,B);
	assign Y = (A&B);
endmodule