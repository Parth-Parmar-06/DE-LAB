module not_1(output Y, input A);
	assign Y = (!A);
endmodule